typedef uvm_sequencer#(wr_tx) write_sqr;
